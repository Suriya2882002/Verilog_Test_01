module and_continous_assignment(input a,input b,output c);
  assign c = a && b;
endmodule
